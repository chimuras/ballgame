module FSM(
	clk,
	xaddr,
	yaddr,
	key_start,
	user1_left,
	user1_right,
	user2_left,
	user2_right,
	score_user1,
	score_user2,
	disp_sel,
	music_en,
	ball_xaddr,
	ball_yaddr,
	user1_xaddr,
	user1_yaddr,
	user2_xaddr,
	user2_yaddr,
	block1_xaddr,
	block1_yaddr,
	block2_xaddr,
	block2_yaddr,
	block3_xaddr,
	block3_yaddr
);

	input			clk;
	input	[9:0] 	xaddr;
	input	[9:0] 	yaddr;
	input			key_start;
	input			user1_left;
	input			user1_right;
	input			user2_left;
	input			user2_right;
	output			disp_sel;
	output			music_en;
	output	[3:0] 	score_user1;
	output	[3:0] 	score_user2;	
	output	[9:0] 	ball_xaddr;
	output	[9:0] 	ball_yaddr;
	output	[9:0] 	user1_xaddr;
	output	[9:0] 	user1_yaddr;
	output	[9:0] 	user2_xaddr;
	output	[9:0] 	user2_yaddr;
	output	[9:0] 	block1_xaddr;
	output	[9:0] 	block1_yaddr;
	output	[9:0] 	block2_xaddr;
	output	[9:0] 	block2_yaddr;
	output	[9:0] 	block3_xaddr;
	output	[9:0] 	block3_yaddr;

	reg		[3:0] 	score_user1=0;
	reg		[3:0] 	score_user2=0;	
	reg		[9:0] 	ball_xaddr=320;
	reg		[9:0] 	ball_yaddr=440;
	reg		[9:0] 	user1_xaddr=320;
	reg		[9:0] 	user1_yaddr=20;
	reg		[9:0] 	user2_xaddr=320;
	reg		[9:0] 	user2_yaddr=460;
	reg		[9:0] 	block1_xaddr=120;
	reg		[9:0] 	block1_yaddr=120;
	reg		[9:0] 	block2_xaddr=320;
	reg		[9:0] 	block2_yaddr=120;
	reg		[9:0] 	block3_xaddr=520;
	reg		[9:0] 	block3_yaddr=120;
		
	parameter    	HIGH_block	= 60;
	parameter    	WIDTH_block = 120;

	parameter    	HIGH_user	= 20;
	parameter    	WIDTH_user	= 120;
	parameter    	STEP  		= 250;
	reg		[39:0]	cnt_div		= 0;
	reg				clk_div		= 0;
	
	reg		[1:0]	ball_dir	= 0;
	reg				ball_move_en= 1;
	reg				ball_reset	= 0;
	
	parameter    	IDLE 	= 3'b001;
	parameter    	RUN		= 3'b010;
	parameter    	OVER	= 3'b100;
	reg	[2:0]		state	= IDLE;
	

	always@(posedge clk)begin
		if(cnt_div<50000000)begin
			cnt_div<=cnt_div+STEP;
			clk_div<=0;
		end
		else begin
			cnt_div<=0;
			clk_div<=1;
		end
	end	
	
	reg	[39:0]		cnt_bolock_move	= 0;
	parameter   	BLOCK_STEP  	= 230;
	reg		[1:0]	block_dir= 0;	
	
	always@(posedge clk)begin
		if(cnt_bolock_move<50000000)begin
			cnt_bolock_move<=cnt_bolock_move+BLOCK_STEP;
		end
		else begin
			cnt_bolock_move<=0;
			case(block_dir)
			0:begin
				if(block1_xaddr<180)begin
					block1_xaddr<=block1_xaddr+1;
					block2_xaddr<=block2_xaddr+1;
					block3_xaddr<=block3_xaddr+1;
					block_dir<=0;
				end
				else begin
					block_dir<=1;
				end	
			end
			1:begin
				if(block1_yaddr>180)begin
					block1_yaddr<=block1_yaddr-1;
					block2_yaddr<=block2_yaddr-1;
					block3_yaddr<=block3_yaddr-1;
					block_dir<=1;
				end
				else begin
					block_dir<=2;
				end					
			end
			2:begin
				if(block1_xaddr>60)begin
					block1_xaddr<=block1_xaddr-1;
					block2_xaddr<=block2_xaddr-1;
					block3_xaddr<=block3_xaddr-1;
					block_dir<=2;
				end
				else begin
					block_dir<=3;
				end				
			end
			3:begin
				if(block1_yaddr<300)begin
					block1_yaddr<=block1_yaddr+1;
					block2_yaddr<=block2_yaddr+1;
					block3_yaddr<=block3_yaddr+1;
					block_dir<=3;
				end
				else begin
					block_dir<=0;
				end			
			end
			endcase								
		end
	end
	
	
	always@(posedge clk)begin
		if(ball_reset==1)begin
			ball_xaddr<=320;
			ball_yaddr<=440;
		end
		else if(ball_move_en==1 && clk_div==1)begin
			case(ball_dir)
			0:begin
				ball_xaddr<=ball_xaddr+1;
				ball_yaddr<=ball_yaddr-1;
			end
			1:begin
				ball_xaddr<=ball_xaddr-1;
				ball_yaddr<=ball_yaddr-1;			
			end
			2:begin
				ball_xaddr<=ball_xaddr-1;
				ball_yaddr<=ball_yaddr+1;			
			end
			3:begin
				ball_xaddr<=ball_xaddr+1;
				ball_yaddr<=ball_yaddr+1;				
			end
			endcase								
		end
	end
	
	always@(posedge clk)begin
		case(ball_dir)
			0:begin
				if(ball_yaddr>=block1_yaddr-HIGH_block/2 && ball_yaddr<=block1_yaddr+HIGH_block/2 && ball_xaddr==block1_xaddr-WIDTH_block/2)
					ball_dir<=1;
				else if(ball_yaddr>=block2_yaddr-HIGH_block/2 && ball_yaddr<=block2_yaddr+HIGH_block/2 && ball_xaddr==block2_xaddr-WIDTH_block/2)
					ball_dir<=1;
				else if(ball_yaddr>=block3_yaddr-HIGH_block/2 && ball_yaddr<=block3_yaddr+HIGH_block/2 && ball_xaddr==block3_xaddr-WIDTH_block/2)
					ball_dir<=1;										
				else if(ball_xaddr==620)
					ball_dir<=1;
				else if(ball_xaddr>=block1_xaddr-WIDTH_block/2 && ball_xaddr<=block1_xaddr+WIDTH_block/2 && ball_yaddr==block1_yaddr+HIGH_block/2)
					ball_dir<=3;
				else if(ball_xaddr>=block2_xaddr-WIDTH_block/2 && ball_xaddr<=block2_xaddr+WIDTH_block/2 && ball_yaddr==block2_yaddr+HIGH_block/2)
					ball_dir<=3;
				else if(ball_xaddr>=block3_xaddr-WIDTH_block/2 && ball_xaddr<=block3_xaddr+WIDTH_block/2 && ball_yaddr==block3_yaddr+HIGH_block/2)
					ball_dir<=3;
				else if(ball_xaddr>=user1_xaddr-WIDTH_user/2 && ball_xaddr<=user1_xaddr+WIDTH_user/2 && ball_yaddr==40)
					ball_dir<=3;															
				else if(ball_yaddr==20)
					ball_dir<=3;
				else
					ball_dir<=0;
			end
			1:begin
				if(ball_yaddr>=block1_yaddr-HIGH_block/2 && ball_yaddr<=block1_yaddr+HIGH_block/2 && ball_xaddr==block1_xaddr+WIDTH_block/2)
					ball_dir<=0;
				else if(ball_yaddr>=block2_yaddr-HIGH_block/2 && ball_yaddr<=block2_yaddr+HIGH_block/2 && ball_xaddr==block2_xaddr+WIDTH_block/2)
					ball_dir<=0;
				else if(ball_yaddr>=block3_yaddr-HIGH_block/2 && ball_yaddr<=block3_yaddr+HIGH_block/2 && ball_xaddr==block3_xaddr+WIDTH_block/2)
					ball_dir<=0;										
				else if(ball_xaddr==20)
					ball_dir<=0;
				else if(ball_xaddr>=block1_xaddr-WIDTH_block/2 && ball_xaddr<=block1_xaddr+WIDTH_block/2 && ball_yaddr==block1_yaddr+HIGH_block/2)
					ball_dir<=2;
				else if(ball_xaddr>=block2_xaddr-WIDTH_block/2 && ball_xaddr<=block2_xaddr+WIDTH_block/2 && ball_yaddr==block2_yaddr+HIGH_block/2)
					ball_dir<=2;
				else if(ball_xaddr>=block3_xaddr-WIDTH_block/2 && ball_xaddr<=block3_xaddr+WIDTH_block/2 && ball_yaddr==block3_yaddr+HIGH_block/2)
					ball_dir<=2;
				else if(ball_xaddr>=user1_xaddr-WIDTH_user/2 && ball_xaddr<=user1_xaddr+WIDTH_user/2 && ball_yaddr==40)
					ball_dir<=2;															
				else if(ball_yaddr==20)
					ball_dir<=2;
				else
					ball_dir<=1;		
			end
			2:begin
				if(ball_yaddr>=block1_yaddr-HIGH_block/2 && ball_yaddr<=block1_yaddr+HIGH_block/2 && ball_xaddr==block1_xaddr+WIDTH_block/2)
					ball_dir<=3;
				else if(ball_yaddr>=block2_yaddr-HIGH_block/2 && ball_yaddr<=block2_yaddr+HIGH_block/2 && ball_xaddr==block2_xaddr+WIDTH_block/2)
					ball_dir<=3;
				else if(ball_yaddr>=block3_yaddr-HIGH_block/2 && ball_yaddr<=block3_yaddr+HIGH_block/2 && ball_xaddr==block3_xaddr+WIDTH_block/2)
					ball_dir<=3;										
				else if(ball_xaddr==20)
					ball_dir<=3;
				else if(ball_xaddr>=block1_xaddr-WIDTH_block/2 && ball_xaddr<=block1_xaddr+WIDTH_block/2 && ball_yaddr==block1_yaddr-HIGH_block/2)
					ball_dir<=1;
				else if(ball_xaddr>=block2_xaddr-WIDTH_block/2 && ball_xaddr<=block2_xaddr+WIDTH_block/2 && ball_yaddr==block2_yaddr-HIGH_block/2)
					ball_dir<=1;
				else if(ball_xaddr>=block3_xaddr-WIDTH_block/2 && ball_xaddr<=block3_xaddr+WIDTH_block/2 && ball_yaddr==block3_yaddr-HIGH_block/2)
					ball_dir<=1;
				else if(ball_xaddr>=user2_xaddr-WIDTH_user/2 && ball_xaddr<=user2_xaddr+WIDTH_user/2 && ball_yaddr==440)
					ball_dir<=1;															
				else if(ball_yaddr==460)
					ball_dir<=1;
				else
					ball_dir<=2;		
			end
			3:begin
				if(ball_yaddr>=block1_yaddr-HIGH_block/2 && ball_yaddr<=block1_yaddr+HIGH_block/2 && ball_xaddr==block1_xaddr-WIDTH_block/2)
					ball_dir<=2;
				else if(ball_yaddr>=block2_yaddr-HIGH_block/2 && ball_yaddr<=block2_yaddr+HIGH_block/2 && ball_xaddr==block2_xaddr-WIDTH_block/2)
					ball_dir<=2;
				else if(ball_yaddr>=block3_yaddr-HIGH_block/2 && ball_yaddr<=block3_yaddr+HIGH_block/2 && ball_xaddr==block3_xaddr-WIDTH_block/2)
					ball_dir<=2;										
				else if(ball_xaddr==620)
					ball_dir<=2;
				else if(ball_xaddr>=block1_xaddr-WIDTH_block/2 && ball_xaddr<=block1_xaddr+WIDTH_block/2 && ball_yaddr==block1_yaddr-HIGH_block/2)
					ball_dir<=0;
				else if(ball_xaddr>=block2_xaddr-WIDTH_block/2 && ball_xaddr<=block2_xaddr+WIDTH_block/2 && ball_yaddr==block2_yaddr-HIGH_block/2)
					ball_dir<=0;
				else if(ball_xaddr>=block3_xaddr-WIDTH_block/2 && ball_xaddr<=block3_xaddr+WIDTH_block/2 && ball_yaddr==block3_yaddr-HIGH_block/2)
					ball_dir<=0;
				else if(ball_xaddr>=user2_xaddr-WIDTH_user/2 && ball_xaddr<=user2_xaddr+WIDTH_user/2 && ball_yaddr==440)
					ball_dir<=0;															
				else if(ball_yaddr==460)
					ball_dir<=0;
				else
					ball_dir<=3;			
			end
		endcase	
	end
	
	always@(posedge clk)begin
		case(state)
			IDLE : begin
				ball_move_en<=0;
				score_user1	<=0;
				score_user2 <=0;
				user1_xaddr <=320;
				user1_yaddr <=20;
				user2_xaddr <=320;
				user2_yaddr <=460;
				ball_reset	<=1;
				if(key_start==1)begin
					state<=RUN;
					ball_move_en<=1;
					ball_reset	<=0;
				end	
				else begin
					state<=IDLE;
				end
			end
			RUN  : begin
				ball_move_en<=1;
				if(ball_reset==0)begin
					if(user1_left==1)begin
						if(user1_xaddr>50)
							user1_xaddr<=user1_xaddr-10;
						else
							user1_xaddr<=50;
					end
					else if(user1_right==1)begin
						if(user1_xaddr<590)
							user1_xaddr<=user1_xaddr+10;
						else
							user1_xaddr<=590;
					end
					if(user2_left==1)begin
						if(user2_xaddr>50)
							user2_xaddr<=user2_xaddr-10;
						else
							user2_xaddr<=50;
					end
					else if(user2_right==1)begin
						if(user2_xaddr<590)
							user2_xaddr<=user2_xaddr+10;
						else
							user2_xaddr<=590;
					end
				end
				if(key_start==1)begin
					ball_reset	<=0;
				end
				if(ball_yaddr<=22)begin
					if(ball_reset==0)begin
						if(score_user1<4)begin
							score_user1<=score_user1+1;
							state<=RUN;
						end
						else begin
							score_user1<=score_user1+1;
							state<=OVER;
						end
					end
					ball_reset	<=1;
					user1_xaddr <=320;
					user1_yaddr <=20;
					user2_xaddr <=320;
					user2_yaddr <=460;					
				end
				else if(ball_yaddr>=458)begin
					if(ball_reset==0)begin
						if(score_user2<4)begin
							score_user2<=score_user2+1;
							state<=RUN;
						end
						else begin
							score_user2<=score_user2+1;
							state<=OVER;
						end
					end
					ball_reset	<=1;
					user1_xaddr <=320;
					user1_yaddr <=20;
					user2_xaddr <=320;
					user2_yaddr <=460;					
				end
				else begin
					state<=RUN;
				end
			end
			OVER : begin
				ball_move_en<=0;
				if(key_start==1)begin
					state<=IDLE;
				end	
				else begin
					state<=OVER;
				end				
			end
		endcase
	end

	assign disp_sel=(state==OVER)? 1'b1 :1'b0;
	assign music_en=(state==RUN)? 1'b1 :1'b0;
//	assign disp_sel=1'b1;

endmodule 						
        